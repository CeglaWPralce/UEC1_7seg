module top (
    // ...
);

// ...

endmodule
